// final_project_soc.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module final_project_soc (
		input  wire        clk_clk,          //        clk.clk
		input  wire [7:0]  keycode_export,   //    keycode.export
		output wire        m1alive_export,   //    m1alive.export
		output wire [11:0] m1posx_export,    //     m1posx.export
		output wire [9:0]  m1posy_export,    //     m1posy.export
		output wire        m2alive_export,   //    m2alive.export
		output wire [11:0] m2posx_export,    //     m2posx.export
		output wire [9:0]  m2posy_export,    //     m2posy.export
		output wire [11:0] mapposx_export,   //    mapposx.export
		output wire        p1_att_export,    //     p1_att.export
		output wire        p1d_export,       //        p1d.export
		output wire [2:0]  p1hp_export,      //       p1hp.export
		output wire [11:0] p1posx_export,    //     p1posx.export
		output wire [9:0]  p1posy_export,    //     p1posy.export
		input  wire        press_export,     //      press.export
		input  wire        reset_reset_n,    //      reset.reset_n
		output wire        rocket_on_export, //  rocket_on.export
		output wire [11:0] rposx_export,     //      rposx.export
		output wire [9:0]  rposy_export,     //      rposy.export
		output wire [4:0]  score_export,     //      score.export
		output wire        sdram_clk_clk,    //  sdram_clk.clk
		output wire [12:0] sdram_wire_addr,  // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,    //           .ba
		output wire        sdram_wire_cas_n, //           .cas_n
		output wire        sdram_wire_cke,   //           .cke
		output wire        sdram_wire_cs_n,  //           .cs_n
		inout  wire [31:0] sdram_wire_dq,    //           .dq
		output wire [3:0]  sdram_wire_dqm,   //           .dqm
		output wire        sdram_wire_ras_n, //           .ras_n
		output wire        sdram_wire_we_n,  //           .we_n
		output wire [1:0]  stage_export,     //      stage.export
		output wire        win_export        //        win.export
	);

	wire         sdram_pll_c0_clk;                                            // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_002:clk, sdram:clk]
	wire  [31:0] nios2_qsys_0_data_master_readdata;                           // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                        // nios2_qsys_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [29:0] nios2_qsys_0_data_master_address;                            // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                         // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                               // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                              // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                          // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [28:0] nios2_qsys_0_instruction_master_address;                     // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                        // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata;     // nios2_qsys_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest;  // nios2_qsys_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_debugaccess -> nios2_qsys_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_address -> nios2_qsys_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_read -> nios2_qsys_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_byteenable -> nios2_qsys_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_write -> nios2_qsys_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_writedata -> nios2_qsys_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;              // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;               // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                  // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                 // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;             // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                       // keyCode:readdata -> mm_interconnect_0:keyCode_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                        // mm_interconnect_0:keyCode_s1_address -> keyCode:address
	wire         mm_interconnect_0_p1posx_s1_chipselect;                      // mm_interconnect_0:p1PosX_s1_chipselect -> p1PosX:chipselect
	wire  [31:0] mm_interconnect_0_p1posx_s1_readdata;                        // p1PosX:readdata -> mm_interconnect_0:p1PosX_s1_readdata
	wire   [1:0] mm_interconnect_0_p1posx_s1_address;                         // mm_interconnect_0:p1PosX_s1_address -> p1PosX:address
	wire         mm_interconnect_0_p1posx_s1_write;                           // mm_interconnect_0:p1PosX_s1_write -> p1PosX:write_n
	wire  [31:0] mm_interconnect_0_p1posx_s1_writedata;                       // mm_interconnect_0:p1PosX_s1_writedata -> p1PosX:writedata
	wire         mm_interconnect_0_p1posy_s1_chipselect;                      // mm_interconnect_0:p1PosY_s1_chipselect -> p1PosY:chipselect
	wire  [31:0] mm_interconnect_0_p1posy_s1_readdata;                        // p1PosY:readdata -> mm_interconnect_0:p1PosY_s1_readdata
	wire   [1:0] mm_interconnect_0_p1posy_s1_address;                         // mm_interconnect_0:p1PosY_s1_address -> p1PosY:address
	wire         mm_interconnect_0_p1posy_s1_write;                           // mm_interconnect_0:p1PosY_s1_write -> p1PosY:write_n
	wire  [31:0] mm_interconnect_0_p1posy_s1_writedata;                       // mm_interconnect_0:p1PosY_s1_writedata -> p1PosY:writedata
	wire         mm_interconnect_0_m1posx_s1_chipselect;                      // mm_interconnect_0:m1PosX_s1_chipselect -> m1PosX:chipselect
	wire  [31:0] mm_interconnect_0_m1posx_s1_readdata;                        // m1PosX:readdata -> mm_interconnect_0:m1PosX_s1_readdata
	wire   [1:0] mm_interconnect_0_m1posx_s1_address;                         // mm_interconnect_0:m1PosX_s1_address -> m1PosX:address
	wire         mm_interconnect_0_m1posx_s1_write;                           // mm_interconnect_0:m1PosX_s1_write -> m1PosX:write_n
	wire  [31:0] mm_interconnect_0_m1posx_s1_writedata;                       // mm_interconnect_0:m1PosX_s1_writedata -> m1PosX:writedata
	wire         mm_interconnect_0_m1posy_s1_chipselect;                      // mm_interconnect_0:m1PosY_s1_chipselect -> m1PosY:chipselect
	wire  [31:0] mm_interconnect_0_m1posy_s1_readdata;                        // m1PosY:readdata -> mm_interconnect_0:m1PosY_s1_readdata
	wire   [1:0] mm_interconnect_0_m1posy_s1_address;                         // mm_interconnect_0:m1PosY_s1_address -> m1PosY:address
	wire         mm_interconnect_0_m1posy_s1_write;                           // mm_interconnect_0:m1PosY_s1_write -> m1PosY:write_n
	wire  [31:0] mm_interconnect_0_m1posy_s1_writedata;                       // mm_interconnect_0:m1PosY_s1_writedata -> m1PosY:writedata
	wire         mm_interconnect_0_p1hp_s1_chipselect;                        // mm_interconnect_0:p1HP_s1_chipselect -> p1HP:chipselect
	wire  [31:0] mm_interconnect_0_p1hp_s1_readdata;                          // p1HP:readdata -> mm_interconnect_0:p1HP_s1_readdata
	wire   [1:0] mm_interconnect_0_p1hp_s1_address;                           // mm_interconnect_0:p1HP_s1_address -> p1HP:address
	wire         mm_interconnect_0_p1hp_s1_write;                             // mm_interconnect_0:p1HP_s1_write -> p1HP:write_n
	wire  [31:0] mm_interconnect_0_p1hp_s1_writedata;                         // mm_interconnect_0:p1HP_s1_writedata -> p1HP:writedata
	wire         mm_interconnect_0_p1_att_s1_chipselect;                      // mm_interconnect_0:p1_Att_s1_chipselect -> p1_Att:chipselect
	wire  [31:0] mm_interconnect_0_p1_att_s1_readdata;                        // p1_Att:readdata -> mm_interconnect_0:p1_Att_s1_readdata
	wire   [1:0] mm_interconnect_0_p1_att_s1_address;                         // mm_interconnect_0:p1_Att_s1_address -> p1_Att:address
	wire         mm_interconnect_0_p1_att_s1_write;                           // mm_interconnect_0:p1_Att_s1_write -> p1_Att:write_n
	wire  [31:0] mm_interconnect_0_p1_att_s1_writedata;                       // mm_interconnect_0:p1_Att_s1_writedata -> p1_Att:writedata
	wire         mm_interconnect_0_p1d_s1_chipselect;                         // mm_interconnect_0:p1D_s1_chipselect -> p1D:chipselect
	wire  [31:0] mm_interconnect_0_p1d_s1_readdata;                           // p1D:readdata -> mm_interconnect_0:p1D_s1_readdata
	wire   [1:0] mm_interconnect_0_p1d_s1_address;                            // mm_interconnect_0:p1D_s1_address -> p1D:address
	wire         mm_interconnect_0_p1d_s1_write;                              // mm_interconnect_0:p1D_s1_write -> p1D:write_n
	wire  [31:0] mm_interconnect_0_p1d_s1_writedata;                          // mm_interconnect_0:p1D_s1_writedata -> p1D:writedata
	wire         mm_interconnect_0_m1alive_s1_chipselect;                     // mm_interconnect_0:m1Alive_s1_chipselect -> m1Alive:chipselect
	wire  [31:0] mm_interconnect_0_m1alive_s1_readdata;                       // m1Alive:readdata -> mm_interconnect_0:m1Alive_s1_readdata
	wire   [1:0] mm_interconnect_0_m1alive_s1_address;                        // mm_interconnect_0:m1Alive_s1_address -> m1Alive:address
	wire         mm_interconnect_0_m1alive_s1_write;                          // mm_interconnect_0:m1Alive_s1_write -> m1Alive:write_n
	wire  [31:0] mm_interconnect_0_m1alive_s1_writedata;                      // mm_interconnect_0:m1Alive_s1_writedata -> m1Alive:writedata
	wire  [31:0] mm_interconnect_0_press_s1_readdata;                         // press:readdata -> mm_interconnect_0:press_s1_readdata
	wire   [1:0] mm_interconnect_0_press_s1_address;                          // mm_interconnect_0:press_s1_address -> press:address
	wire         mm_interconnect_0_m2posx_s1_chipselect;                      // mm_interconnect_0:m2PosX_s1_chipselect -> m2PosX:chipselect
	wire  [31:0] mm_interconnect_0_m2posx_s1_readdata;                        // m2PosX:readdata -> mm_interconnect_0:m2PosX_s1_readdata
	wire   [1:0] mm_interconnect_0_m2posx_s1_address;                         // mm_interconnect_0:m2PosX_s1_address -> m2PosX:address
	wire         mm_interconnect_0_m2posx_s1_write;                           // mm_interconnect_0:m2PosX_s1_write -> m2PosX:write_n
	wire  [31:0] mm_interconnect_0_m2posx_s1_writedata;                       // mm_interconnect_0:m2PosX_s1_writedata -> m2PosX:writedata
	wire         mm_interconnect_0_m2posy_s1_chipselect;                      // mm_interconnect_0:m2PosY_s1_chipselect -> m2PosY:chipselect
	wire  [31:0] mm_interconnect_0_m2posy_s1_readdata;                        // m2PosY:readdata -> mm_interconnect_0:m2PosY_s1_readdata
	wire   [1:0] mm_interconnect_0_m2posy_s1_address;                         // mm_interconnect_0:m2PosY_s1_address -> m2PosY:address
	wire         mm_interconnect_0_m2posy_s1_write;                           // mm_interconnect_0:m2PosY_s1_write -> m2PosY:write_n
	wire  [31:0] mm_interconnect_0_m2posy_s1_writedata;                       // mm_interconnect_0:m2PosY_s1_writedata -> m2PosY:writedata
	wire         mm_interconnect_0_m2alive_s1_chipselect;                     // mm_interconnect_0:m2Alive_s1_chipselect -> m2Alive:chipselect
	wire  [31:0] mm_interconnect_0_m2alive_s1_readdata;                       // m2Alive:readdata -> mm_interconnect_0:m2Alive_s1_readdata
	wire   [1:0] mm_interconnect_0_m2alive_s1_address;                        // mm_interconnect_0:m2Alive_s1_address -> m2Alive:address
	wire         mm_interconnect_0_m2alive_s1_write;                          // mm_interconnect_0:m2Alive_s1_write -> m2Alive:write_n
	wire  [31:0] mm_interconnect_0_m2alive_s1_writedata;                      // mm_interconnect_0:m2Alive_s1_writedata -> m2Alive:writedata
	wire         mm_interconnect_0_mapposx_s1_chipselect;                     // mm_interconnect_0:mapPosX_s1_chipselect -> mapPosX:chipselect
	wire  [31:0] mm_interconnect_0_mapposx_s1_readdata;                       // mapPosX:readdata -> mm_interconnect_0:mapPosX_s1_readdata
	wire   [1:0] mm_interconnect_0_mapposx_s1_address;                        // mm_interconnect_0:mapPosX_s1_address -> mapPosX:address
	wire         mm_interconnect_0_mapposx_s1_write;                          // mm_interconnect_0:mapPosX_s1_write -> mapPosX:write_n
	wire  [31:0] mm_interconnect_0_mapposx_s1_writedata;                      // mm_interconnect_0:mapPosX_s1_writedata -> mapPosX:writedata
	wire         mm_interconnect_0_rposx_s1_chipselect;                       // mm_interconnect_0:rPosX_s1_chipselect -> rPosX:chipselect
	wire  [31:0] mm_interconnect_0_rposx_s1_readdata;                         // rPosX:readdata -> mm_interconnect_0:rPosX_s1_readdata
	wire   [1:0] mm_interconnect_0_rposx_s1_address;                          // mm_interconnect_0:rPosX_s1_address -> rPosX:address
	wire         mm_interconnect_0_rposx_s1_write;                            // mm_interconnect_0:rPosX_s1_write -> rPosX:write_n
	wire  [31:0] mm_interconnect_0_rposx_s1_writedata;                        // mm_interconnect_0:rPosX_s1_writedata -> rPosX:writedata
	wire         mm_interconnect_0_rposy_s1_chipselect;                       // mm_interconnect_0:rPosY_s1_chipselect -> rPosY:chipselect
	wire  [31:0] mm_interconnect_0_rposy_s1_readdata;                         // rPosY:readdata -> mm_interconnect_0:rPosY_s1_readdata
	wire   [1:0] mm_interconnect_0_rposy_s1_address;                          // mm_interconnect_0:rPosY_s1_address -> rPosY:address
	wire         mm_interconnect_0_rposy_s1_write;                            // mm_interconnect_0:rPosY_s1_write -> rPosY:write_n
	wire  [31:0] mm_interconnect_0_rposy_s1_writedata;                        // mm_interconnect_0:rPosY_s1_writedata -> rPosY:writedata
	wire         mm_interconnect_0_rocket_on_s1_chipselect;                   // mm_interconnect_0:rocket_on_s1_chipselect -> rocket_on:chipselect
	wire  [31:0] mm_interconnect_0_rocket_on_s1_readdata;                     // rocket_on:readdata -> mm_interconnect_0:rocket_on_s1_readdata
	wire   [1:0] mm_interconnect_0_rocket_on_s1_address;                      // mm_interconnect_0:rocket_on_s1_address -> rocket_on:address
	wire         mm_interconnect_0_rocket_on_s1_write;                        // mm_interconnect_0:rocket_on_s1_write -> rocket_on:write_n
	wire  [31:0] mm_interconnect_0_rocket_on_s1_writedata;                    // mm_interconnect_0:rocket_on_s1_writedata -> rocket_on:writedata
	wire         mm_interconnect_0_score_s1_chipselect;                       // mm_interconnect_0:Score_s1_chipselect -> Score:chipselect
	wire  [31:0] mm_interconnect_0_score_s1_readdata;                         // Score:readdata -> mm_interconnect_0:Score_s1_readdata
	wire   [1:0] mm_interconnect_0_score_s1_address;                          // mm_interconnect_0:Score_s1_address -> Score:address
	wire         mm_interconnect_0_score_s1_write;                            // mm_interconnect_0:Score_s1_write -> Score:write_n
	wire  [31:0] mm_interconnect_0_score_s1_writedata;                        // mm_interconnect_0:Score_s1_writedata -> Score:writedata
	wire         mm_interconnect_0_stage_s1_chipselect;                       // mm_interconnect_0:stage_s1_chipselect -> stage:chipselect
	wire  [31:0] mm_interconnect_0_stage_s1_readdata;                         // stage:readdata -> mm_interconnect_0:stage_s1_readdata
	wire   [1:0] mm_interconnect_0_stage_s1_address;                          // mm_interconnect_0:stage_s1_address -> stage:address
	wire         mm_interconnect_0_stage_s1_write;                            // mm_interconnect_0:stage_s1_write -> stage:write_n
	wire  [31:0] mm_interconnect_0_stage_s1_writedata;                        // mm_interconnect_0:stage_s1_writedata -> stage:writedata
	wire         mm_interconnect_0_win_s1_chipselect;                         // mm_interconnect_0:win_s1_chipselect -> win:chipselect
	wire  [31:0] mm_interconnect_0_win_s1_readdata;                           // win:readdata -> mm_interconnect_0:win_s1_readdata
	wire   [1:0] mm_interconnect_0_win_s1_address;                            // mm_interconnect_0:win_s1_address -> win:address
	wire         mm_interconnect_0_win_s1_write;                              // mm_interconnect_0:win_s1_write -> win:write_n
	wire  [31:0] mm_interconnect_0_win_s1_writedata;                          // mm_interconnect_0:win_s1_writedata -> win:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_qsys_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Score:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, keyCode:reset_n, m1Alive:reset_n, m1PosX:reset_n, m1PosY:reset_n, m2Alive:reset_n, m2PosX:reset_n, m2PosY:reset_n, mapPosX:reset_n, mm_interconnect_0:nios2_qsys_0_reset_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, p1D:reset_n, p1HP:reset_n, p1PosX:reset_n, p1PosY:reset_n, p1_Att:reset_n, press:reset_n, rPosX:reset_n, rPosY:reset_n, rocket_on:reset_n, rst_translator:in_reset, stage:reset_n, win:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_qsys_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_debug_reset_request_reset;                      // nios2_qsys_0:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:sysid_qsys_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator_001:in_reset, sdram_pll:reset, sysid_qsys_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [onchip_memory2_0:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	final_project_soc_Score score (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_score_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_score_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_score_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_score_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_score_s1_readdata),   //                    .readdata
		.out_port   (score_export)                           // external_connection.export
	);

	final_project_soc_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	final_project_soc_keyCode keycode (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_keycode_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_keycode_s1_readdata), //                    .readdata
		.in_port  (keycode_export)                         // external_connection.export
	);

	final_project_soc_m1Alive m1alive (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_m1alive_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_m1alive_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_m1alive_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_m1alive_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_m1alive_s1_readdata),   //                    .readdata
		.out_port   (m1alive_export)                           // external_connection.export
	);

	final_project_soc_m1PosX m1posx (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_m1posx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_m1posx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_m1posx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_m1posx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_m1posx_s1_readdata),   //                    .readdata
		.out_port   (m1posx_export)                           // external_connection.export
	);

	final_project_soc_m1PosY m1posy (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_m1posy_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_m1posy_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_m1posy_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_m1posy_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_m1posy_s1_readdata),   //                    .readdata
		.out_port   (m1posy_export)                           // external_connection.export
	);

	final_project_soc_m1Alive m2alive (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_m2alive_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_m2alive_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_m2alive_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_m2alive_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_m2alive_s1_readdata),   //                    .readdata
		.out_port   (m2alive_export)                           // external_connection.export
	);

	final_project_soc_m1PosX m2posx (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_m2posx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_m2posx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_m2posx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_m2posx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_m2posx_s1_readdata),   //                    .readdata
		.out_port   (m2posx_export)                           // external_connection.export
	);

	final_project_soc_m1PosY m2posy (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_m2posy_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_m2posy_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_m2posy_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_m2posy_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_m2posy_s1_readdata),   //                    .readdata
		.out_port   (m2posy_export)                           // external_connection.export
	);

	final_project_soc_m1PosX mapposx (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_mapposx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mapposx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mapposx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mapposx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mapposx_s1_readdata),   //                    .readdata
		.out_port   (mapposx_export)                           // external_connection.export
	);

	final_project_soc_nios2_qsys_0 nios2_qsys_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_qsys_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_qsys_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_qsys_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	final_project_soc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)            //       .reset_req
	);

	final_project_soc_m1Alive p1d (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_p1d_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_p1d_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_p1d_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_p1d_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_p1d_s1_readdata),   //                    .readdata
		.out_port   (p1d_export)                           // external_connection.export
	);

	final_project_soc_p1HP p1hp (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_p1hp_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_p1hp_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_p1hp_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_p1hp_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_p1hp_s1_readdata),   //                    .readdata
		.out_port   (p1hp_export)                           // external_connection.export
	);

	final_project_soc_m1PosX p1posx (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_p1posx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_p1posx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_p1posx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_p1posx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_p1posx_s1_readdata),   //                    .readdata
		.out_port   (p1posx_export)                           // external_connection.export
	);

	final_project_soc_m1PosY p1posy (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_p1posy_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_p1posy_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_p1posy_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_p1posy_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_p1posy_s1_readdata),   //                    .readdata
		.out_port   (p1posy_export)                           // external_connection.export
	);

	final_project_soc_m1Alive p1_att (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_p1_att_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_p1_att_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_p1_att_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_p1_att_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_p1_att_s1_readdata),   //                    .readdata
		.out_port   (p1_att_export)                           // external_connection.export
	);

	final_project_soc_press press (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_press_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_press_s1_readdata), //                    .readdata
		.in_port  (press_export)                         // external_connection.export
	);

	final_project_soc_m1PosX rposx (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_rposx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rposx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rposx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rposx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rposx_s1_readdata),   //                    .readdata
		.out_port   (rposx_export)                           // external_connection.export
	);

	final_project_soc_m1PosY rposy (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_rposy_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rposy_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rposy_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rposy_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rposy_s1_readdata),   //                    .readdata
		.out_port   (rposy_export)                           // external_connection.export
	);

	final_project_soc_m1Alive rocket_on (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_rocket_on_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rocket_on_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rocket_on_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rocket_on_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rocket_on_s1_readdata),   //                    .readdata
		.out_port   (rocket_on_export)                           // external_connection.export
	);

	final_project_soc_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	final_project_soc_sdram_pll sdram_pll (
		.clk       (clk_clk),                                         //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),              // inclk_interface_reset.reset
		.read      (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0        (sdram_pll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                                   //                    c1.clk
		.areset    (),                                                //        areset_conduit.export
		.locked    (),                                                //        locked_conduit.export
		.phasedone ()                                                 //     phasedone_conduit.export
	);

	final_project_soc_stage stage (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_stage_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_stage_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_stage_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_stage_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_stage_s1_readdata),   //                    .readdata
		.out_port   (stage_export)                           // external_connection.export
	);

	final_project_soc_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	final_project_soc_m1Alive win (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_win_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_win_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_win_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_win_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_win_s1_readdata),   //                    .readdata
		.out_port   (win_export)                           // external_connection.export
	);

	final_project_soc_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.sdram_pll_c0_clk                               (sdram_pll_c0_clk),                                            //                             sdram_pll_c0.clk
		.nios2_qsys_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_qsys_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset        (rst_controller_002_reset_out_reset),                          //        sdram_reset_reset_bridge_in_reset.reset
		.sysid_qsys_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // sysid_qsys_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address               (nios2_qsys_0_data_master_address),                            //                 nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest           (nios2_qsys_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_qsys_0_data_master_byteenable            (nios2_qsys_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_qsys_0_data_master_read                  (nios2_qsys_0_data_master_read),                               //                                         .read
		.nios2_qsys_0_data_master_readdata              (nios2_qsys_0_data_master_readdata),                           //                                         .readdata
		.nios2_qsys_0_data_master_write                 (nios2_qsys_0_data_master_write),                              //                                         .write
		.nios2_qsys_0_data_master_writedata             (nios2_qsys_0_data_master_writedata),                          //                                         .writedata
		.nios2_qsys_0_data_master_debugaccess           (nios2_qsys_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_qsys_0_instruction_master_address        (nios2_qsys_0_instruction_master_address),                     //          nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest    (nios2_qsys_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_qsys_0_instruction_master_read           (nios2_qsys_0_instruction_master_read),                        //                                         .read
		.nios2_qsys_0_instruction_master_readdata       (nios2_qsys_0_instruction_master_readdata),                    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.keyCode_s1_address                             (mm_interconnect_0_keycode_s1_address),                        //                               keyCode_s1.address
		.keyCode_s1_readdata                            (mm_interconnect_0_keycode_s1_readdata),                       //                                         .readdata
		.m1Alive_s1_address                             (mm_interconnect_0_m1alive_s1_address),                        //                               m1Alive_s1.address
		.m1Alive_s1_write                               (mm_interconnect_0_m1alive_s1_write),                          //                                         .write
		.m1Alive_s1_readdata                            (mm_interconnect_0_m1alive_s1_readdata),                       //                                         .readdata
		.m1Alive_s1_writedata                           (mm_interconnect_0_m1alive_s1_writedata),                      //                                         .writedata
		.m1Alive_s1_chipselect                          (mm_interconnect_0_m1alive_s1_chipselect),                     //                                         .chipselect
		.m1PosX_s1_address                              (mm_interconnect_0_m1posx_s1_address),                         //                                m1PosX_s1.address
		.m1PosX_s1_write                                (mm_interconnect_0_m1posx_s1_write),                           //                                         .write
		.m1PosX_s1_readdata                             (mm_interconnect_0_m1posx_s1_readdata),                        //                                         .readdata
		.m1PosX_s1_writedata                            (mm_interconnect_0_m1posx_s1_writedata),                       //                                         .writedata
		.m1PosX_s1_chipselect                           (mm_interconnect_0_m1posx_s1_chipselect),                      //                                         .chipselect
		.m1PosY_s1_address                              (mm_interconnect_0_m1posy_s1_address),                         //                                m1PosY_s1.address
		.m1PosY_s1_write                                (mm_interconnect_0_m1posy_s1_write),                           //                                         .write
		.m1PosY_s1_readdata                             (mm_interconnect_0_m1posy_s1_readdata),                        //                                         .readdata
		.m1PosY_s1_writedata                            (mm_interconnect_0_m1posy_s1_writedata),                       //                                         .writedata
		.m1PosY_s1_chipselect                           (mm_interconnect_0_m1posy_s1_chipselect),                      //                                         .chipselect
		.m2Alive_s1_address                             (mm_interconnect_0_m2alive_s1_address),                        //                               m2Alive_s1.address
		.m2Alive_s1_write                               (mm_interconnect_0_m2alive_s1_write),                          //                                         .write
		.m2Alive_s1_readdata                            (mm_interconnect_0_m2alive_s1_readdata),                       //                                         .readdata
		.m2Alive_s1_writedata                           (mm_interconnect_0_m2alive_s1_writedata),                      //                                         .writedata
		.m2Alive_s1_chipselect                          (mm_interconnect_0_m2alive_s1_chipselect),                     //                                         .chipselect
		.m2PosX_s1_address                              (mm_interconnect_0_m2posx_s1_address),                         //                                m2PosX_s1.address
		.m2PosX_s1_write                                (mm_interconnect_0_m2posx_s1_write),                           //                                         .write
		.m2PosX_s1_readdata                             (mm_interconnect_0_m2posx_s1_readdata),                        //                                         .readdata
		.m2PosX_s1_writedata                            (mm_interconnect_0_m2posx_s1_writedata),                       //                                         .writedata
		.m2PosX_s1_chipselect                           (mm_interconnect_0_m2posx_s1_chipselect),                      //                                         .chipselect
		.m2PosY_s1_address                              (mm_interconnect_0_m2posy_s1_address),                         //                                m2PosY_s1.address
		.m2PosY_s1_write                                (mm_interconnect_0_m2posy_s1_write),                           //                                         .write
		.m2PosY_s1_readdata                             (mm_interconnect_0_m2posy_s1_readdata),                        //                                         .readdata
		.m2PosY_s1_writedata                            (mm_interconnect_0_m2posy_s1_writedata),                       //                                         .writedata
		.m2PosY_s1_chipselect                           (mm_interconnect_0_m2posy_s1_chipselect),                      //                                         .chipselect
		.mapPosX_s1_address                             (mm_interconnect_0_mapposx_s1_address),                        //                               mapPosX_s1.address
		.mapPosX_s1_write                               (mm_interconnect_0_mapposx_s1_write),                          //                                         .write
		.mapPosX_s1_readdata                            (mm_interconnect_0_mapposx_s1_readdata),                       //                                         .readdata
		.mapPosX_s1_writedata                           (mm_interconnect_0_mapposx_s1_writedata),                      //                                         .writedata
		.mapPosX_s1_chipselect                          (mm_interconnect_0_mapposx_s1_chipselect),                     //                                         .chipselect
		.nios2_qsys_0_debug_mem_slave_address           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),      //             nios2_qsys_0_debug_mem_slave.address
		.nios2_qsys_0_debug_mem_slave_write             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),        //                                         .write
		.nios2_qsys_0_debug_mem_slave_read              (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),         //                                         .read
		.nios2_qsys_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_qsys_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_qsys_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_qsys_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_qsys_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.p1_Att_s1_address                              (mm_interconnect_0_p1_att_s1_address),                         //                                p1_Att_s1.address
		.p1_Att_s1_write                                (mm_interconnect_0_p1_att_s1_write),                           //                                         .write
		.p1_Att_s1_readdata                             (mm_interconnect_0_p1_att_s1_readdata),                        //                                         .readdata
		.p1_Att_s1_writedata                            (mm_interconnect_0_p1_att_s1_writedata),                       //                                         .writedata
		.p1_Att_s1_chipselect                           (mm_interconnect_0_p1_att_s1_chipselect),                      //                                         .chipselect
		.p1D_s1_address                                 (mm_interconnect_0_p1d_s1_address),                            //                                   p1D_s1.address
		.p1D_s1_write                                   (mm_interconnect_0_p1d_s1_write),                              //                                         .write
		.p1D_s1_readdata                                (mm_interconnect_0_p1d_s1_readdata),                           //                                         .readdata
		.p1D_s1_writedata                               (mm_interconnect_0_p1d_s1_writedata),                          //                                         .writedata
		.p1D_s1_chipselect                              (mm_interconnect_0_p1d_s1_chipselect),                         //                                         .chipselect
		.p1HP_s1_address                                (mm_interconnect_0_p1hp_s1_address),                           //                                  p1HP_s1.address
		.p1HP_s1_write                                  (mm_interconnect_0_p1hp_s1_write),                             //                                         .write
		.p1HP_s1_readdata                               (mm_interconnect_0_p1hp_s1_readdata),                          //                                         .readdata
		.p1HP_s1_writedata                              (mm_interconnect_0_p1hp_s1_writedata),                         //                                         .writedata
		.p1HP_s1_chipselect                             (mm_interconnect_0_p1hp_s1_chipselect),                        //                                         .chipselect
		.p1PosX_s1_address                              (mm_interconnect_0_p1posx_s1_address),                         //                                p1PosX_s1.address
		.p1PosX_s1_write                                (mm_interconnect_0_p1posx_s1_write),                           //                                         .write
		.p1PosX_s1_readdata                             (mm_interconnect_0_p1posx_s1_readdata),                        //                                         .readdata
		.p1PosX_s1_writedata                            (mm_interconnect_0_p1posx_s1_writedata),                       //                                         .writedata
		.p1PosX_s1_chipselect                           (mm_interconnect_0_p1posx_s1_chipselect),                      //                                         .chipselect
		.p1PosY_s1_address                              (mm_interconnect_0_p1posy_s1_address),                         //                                p1PosY_s1.address
		.p1PosY_s1_write                                (mm_interconnect_0_p1posy_s1_write),                           //                                         .write
		.p1PosY_s1_readdata                             (mm_interconnect_0_p1posy_s1_readdata),                        //                                         .readdata
		.p1PosY_s1_writedata                            (mm_interconnect_0_p1posy_s1_writedata),                       //                                         .writedata
		.p1PosY_s1_chipselect                           (mm_interconnect_0_p1posy_s1_chipselect),                      //                                         .chipselect
		.press_s1_address                               (mm_interconnect_0_press_s1_address),                          //                                 press_s1.address
		.press_s1_readdata                              (mm_interconnect_0_press_s1_readdata),                         //                                         .readdata
		.rocket_on_s1_address                           (mm_interconnect_0_rocket_on_s1_address),                      //                             rocket_on_s1.address
		.rocket_on_s1_write                             (mm_interconnect_0_rocket_on_s1_write),                        //                                         .write
		.rocket_on_s1_readdata                          (mm_interconnect_0_rocket_on_s1_readdata),                     //                                         .readdata
		.rocket_on_s1_writedata                         (mm_interconnect_0_rocket_on_s1_writedata),                    //                                         .writedata
		.rocket_on_s1_chipselect                        (mm_interconnect_0_rocket_on_s1_chipselect),                   //                                         .chipselect
		.rPosX_s1_address                               (mm_interconnect_0_rposx_s1_address),                          //                                 rPosX_s1.address
		.rPosX_s1_write                                 (mm_interconnect_0_rposx_s1_write),                            //                                         .write
		.rPosX_s1_readdata                              (mm_interconnect_0_rposx_s1_readdata),                         //                                         .readdata
		.rPosX_s1_writedata                             (mm_interconnect_0_rposx_s1_writedata),                        //                                         .writedata
		.rPosX_s1_chipselect                            (mm_interconnect_0_rposx_s1_chipselect),                       //                                         .chipselect
		.rPosY_s1_address                               (mm_interconnect_0_rposy_s1_address),                          //                                 rPosY_s1.address
		.rPosY_s1_write                                 (mm_interconnect_0_rposy_s1_write),                            //                                         .write
		.rPosY_s1_readdata                              (mm_interconnect_0_rposy_s1_readdata),                         //                                         .readdata
		.rPosY_s1_writedata                             (mm_interconnect_0_rposy_s1_writedata),                        //                                         .writedata
		.rPosY_s1_chipselect                            (mm_interconnect_0_rposy_s1_chipselect),                       //                                         .chipselect
		.Score_s1_address                               (mm_interconnect_0_score_s1_address),                          //                                 Score_s1.address
		.Score_s1_write                                 (mm_interconnect_0_score_s1_write),                            //                                         .write
		.Score_s1_readdata                              (mm_interconnect_0_score_s1_readdata),                         //                                         .readdata
		.Score_s1_writedata                             (mm_interconnect_0_score_s1_writedata),                        //                                         .writedata
		.Score_s1_chipselect                            (mm_interconnect_0_score_s1_chipselect),                       //                                         .chipselect
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                          //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                            //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                             //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                         //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                        //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                       //                                         .chipselect
		.sdram_pll_pll_slave_address                    (mm_interconnect_0_sdram_pll_pll_slave_address),               //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                      (mm_interconnect_0_sdram_pll_pll_slave_write),                 //                                         .write
		.sdram_pll_pll_slave_read                       (mm_interconnect_0_sdram_pll_pll_slave_read),                  //                                         .read
		.sdram_pll_pll_slave_readdata                   (mm_interconnect_0_sdram_pll_pll_slave_readdata),              //                                         .readdata
		.sdram_pll_pll_slave_writedata                  (mm_interconnect_0_sdram_pll_pll_slave_writedata),             //                                         .writedata
		.stage_s1_address                               (mm_interconnect_0_stage_s1_address),                          //                                 stage_s1.address
		.stage_s1_write                                 (mm_interconnect_0_stage_s1_write),                            //                                         .write
		.stage_s1_readdata                              (mm_interconnect_0_stage_s1_readdata),                         //                                         .readdata
		.stage_s1_writedata                             (mm_interconnect_0_stage_s1_writedata),                        //                                         .writedata
		.stage_s1_chipselect                            (mm_interconnect_0_stage_s1_chipselect),                       //                                         .chipselect
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                         .readdata
		.win_s1_address                                 (mm_interconnect_0_win_s1_address),                            //                                   win_s1.address
		.win_s1_write                                   (mm_interconnect_0_win_s1_write),                              //                                         .write
		.win_s1_readdata                                (mm_interconnect_0_win_s1_readdata),                           //                                         .readdata
		.win_s1_writedata                               (mm_interconnect_0_win_s1_writedata),                          //                                         .writedata
		.win_s1_chipselect                              (mm_interconnect_0_win_s1_chipselect)                          //                                         .chipselect
	);

	final_project_soc_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_qsys_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sdram_pll_c0_clk),                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
